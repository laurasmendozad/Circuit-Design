** sch_path: /home/laura/Documents/Circuit Design/Inverter/xschem/inverter_tb.sch
**.subckt inverter_tb out in
*.opin out
*.opin in
*.subckt inverter in vss vdd out
x1 in GND net1 out inverter
V1 in GND PWL(0 0 20n 0 900n 1.8)
V2 net1 GND 1.8
**** begin user architecture code

.lib /home/laura/Documents/ic_design/OpenPDK/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt


.control
tran 1n 1u
plot V(in) V(out)
.endc

**** end user architecture code
**.ends

.include inverter.spice

.GLOBAL GND
.end
